//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company : AGH University of Krakow
// Create Date : 25.08.2024
// Designers Name : Tomasz Ochamenk & Jan PAnek
// Module Name : game_logic
// Project Name : 
// Target Devices : BASYS3
// 
// Description : logika gry, sterowanie 
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module game_logic 
(
    input logic clk,
    input logic rst,
    input logic [1:0] game_board [0:9][0:9],


);


endmodule